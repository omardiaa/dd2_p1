`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//For testing 
//////////////////////////////////////////////////////////////////////////////////

module full_adder #(parameter x=0) (input A,B,cin, output sum, cout);
   
  assign {cout, sum}= A+B+cin;
endmodule
