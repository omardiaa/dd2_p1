`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//For testing 
//////////////////////////////////////////////////////////////////////////////////

module multi_bit_adder  (input[5:0] A,B, input cin, output sum, cout);
   
  assign {cout, sum}= A+B+cin;
endmodule
