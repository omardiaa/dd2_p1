`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//For testing 
//////////////////////////////////////////////////////////////////////////////////

module full_adder #(parameter x=0) (
   input  [5:0] a,
   input  b,
   input  cin,
   output sum,
   output cout
);

   assign {cout,sum} = a+b+cin;
  
endmodule

